--excersize 2 (using structural modeling)

library IEEE;
use IEEE.std_logic_1164.all;


